library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Optional is
  port(clk : in std_logic;
	   en : in std_logic;
	   sel : in std_logic;
	   seed : in std_logic_vector(63 downto 0);
       result : out std_logic_vector(4 downto 0)
  );
end Optional;

architecture behavior of Optional is
  component RNG is
    port(seed : in std_logic_vector(63 downto 0);
         clk, sel : in std_logic;
         rng_out : out std_logic_vector(63 downto 0)
    );
  end component;

  signal rng_output : std_logic_vector(63 downto 0);
  signal mod_output : std_logic_vector(4 downto 0);
  
  -- D Flip-Flop
  signal register_q : std_logic_vector(4 downto 0);

begin
  -- Instantiate the RNG
  RNG_inst : RNG port map(seed => seed,
                           clk => clk,
                           sel => sel,
                           rng_out => rng_output);
  
  -- Modulo-by-21 circuit
  process(clk)
    variable dec_value : integer;
  begin
	if rising_edge(clk) then
		dec_value := to_integer(unsigned(rng_output));

		mod_output <= std_logic_vector(to_unsigned(dec_value mod 21, mod_output'length));
	end if;
  end process;

  -- Register
  process (clk)
  begin
    if rising_edge(clk) then
      if en = '1' then
        register_q <= mod_output;
      end if;
    end if;
  end process;


  -- Output the lottery number
  result <= register_q;

end behavior;